magic
tech sky130A
magscale 1 2
timestamp 1654774612
<< obsli1 >>
rect 1104 2159 178848 117521
<< obsm1 >>
rect 1104 2128 178848 117904
<< metal2 >>
rect 2318 119200 2374 120000
rect 7010 119200 7066 120000
rect 11794 119200 11850 120000
rect 16486 119200 16542 120000
rect 21270 119200 21326 120000
rect 25962 119200 26018 120000
rect 30746 119200 30802 120000
rect 35438 119200 35494 120000
rect 40222 119200 40278 120000
rect 44914 119200 44970 120000
rect 49698 119200 49754 120000
rect 54390 119200 54446 120000
rect 59174 119200 59230 120000
rect 63866 119200 63922 120000
rect 68650 119200 68706 120000
rect 73342 119200 73398 120000
rect 78126 119200 78182 120000
rect 82818 119200 82874 120000
rect 87602 119200 87658 120000
rect 92294 119200 92350 120000
rect 97078 119200 97134 120000
rect 101770 119200 101826 120000
rect 106554 119200 106610 120000
rect 111246 119200 111302 120000
rect 116030 119200 116086 120000
rect 120722 119200 120778 120000
rect 125506 119200 125562 120000
rect 130198 119200 130254 120000
rect 134982 119200 135038 120000
rect 139674 119200 139730 120000
rect 144458 119200 144514 120000
rect 149150 119200 149206 120000
rect 153934 119200 153990 120000
rect 158626 119200 158682 120000
rect 163410 119200 163466 120000
rect 168102 119200 168158 120000
rect 172886 119200 172942 120000
rect 177578 119200 177634 120000
rect 3698 0 3754 800
rect 11150 0 11206 800
rect 18694 0 18750 800
rect 26146 0 26202 800
rect 33690 0 33746 800
rect 41142 0 41198 800
rect 48686 0 48742 800
rect 56138 0 56194 800
rect 63682 0 63738 800
rect 71134 0 71190 800
rect 78678 0 78734 800
rect 86130 0 86186 800
rect 93674 0 93730 800
rect 101218 0 101274 800
rect 108670 0 108726 800
rect 116214 0 116270 800
rect 123666 0 123722 800
rect 131210 0 131266 800
rect 138662 0 138718 800
rect 146206 0 146262 800
rect 153658 0 153714 800
rect 161202 0 161258 800
rect 168654 0 168710 800
rect 176198 0 176254 800
<< obsm2 >>
rect 1398 119144 2262 119354
rect 2430 119144 6954 119354
rect 7122 119144 11738 119354
rect 11906 119144 16430 119354
rect 16598 119144 21214 119354
rect 21382 119144 25906 119354
rect 26074 119144 30690 119354
rect 30858 119144 35382 119354
rect 35550 119144 40166 119354
rect 40334 119144 44858 119354
rect 45026 119144 49642 119354
rect 49810 119144 54334 119354
rect 54502 119144 59118 119354
rect 59286 119144 63810 119354
rect 63978 119144 68594 119354
rect 68762 119144 73286 119354
rect 73454 119144 78070 119354
rect 78238 119144 82762 119354
rect 82930 119144 87546 119354
rect 87714 119144 92238 119354
rect 92406 119144 97022 119354
rect 97190 119144 101714 119354
rect 101882 119144 106498 119354
rect 106666 119144 111190 119354
rect 111358 119144 115974 119354
rect 116142 119144 120666 119354
rect 120834 119144 125450 119354
rect 125618 119144 130142 119354
rect 130310 119144 134926 119354
rect 135094 119144 139618 119354
rect 139786 119144 144402 119354
rect 144570 119144 149094 119354
rect 149262 119144 153878 119354
rect 154046 119144 158570 119354
rect 158738 119144 163354 119354
rect 163522 119144 168046 119354
rect 168214 119144 172830 119354
rect 172998 119144 177522 119354
rect 177690 119144 178186 119354
rect 1398 856 178186 119144
rect 1398 800 3642 856
rect 3810 800 11094 856
rect 11262 800 18638 856
rect 18806 800 26090 856
rect 26258 800 33634 856
rect 33802 800 41086 856
rect 41254 800 48630 856
rect 48798 800 56082 856
rect 56250 800 63626 856
rect 63794 800 71078 856
rect 71246 800 78622 856
rect 78790 800 86074 856
rect 86242 800 93618 856
rect 93786 800 101162 856
rect 101330 800 108614 856
rect 108782 800 116158 856
rect 116326 800 123610 856
rect 123778 800 131154 856
rect 131322 800 138606 856
rect 138774 800 146150 856
rect 146318 800 153602 856
rect 153770 800 161146 856
rect 161314 800 168598 856
rect 168766 800 176142 856
rect 176310 800 178186 856
<< metal3 >>
rect 179200 117648 180000 117768
rect 0 117376 800 117496
rect 179200 113160 180000 113280
rect 0 112344 800 112464
rect 179200 108808 180000 108928
rect 0 107312 800 107432
rect 179200 104320 180000 104440
rect 0 102416 800 102536
rect 179200 99832 180000 99952
rect 0 97384 800 97504
rect 179200 95480 180000 95600
rect 0 92352 800 92472
rect 179200 90992 180000 91112
rect 0 87320 800 87440
rect 179200 86504 180000 86624
rect 0 82424 800 82544
rect 179200 82152 180000 82272
rect 179200 77664 180000 77784
rect 0 77392 800 77512
rect 179200 73176 180000 73296
rect 0 72360 800 72480
rect 179200 68824 180000 68944
rect 0 67328 800 67448
rect 179200 64336 180000 64456
rect 0 62432 800 62552
rect 179200 59848 180000 59968
rect 0 57400 800 57520
rect 179200 55496 180000 55616
rect 0 52368 800 52488
rect 179200 51008 180000 51128
rect 0 47336 800 47456
rect 179200 46520 180000 46640
rect 0 42440 800 42560
rect 179200 42168 180000 42288
rect 179200 37680 180000 37800
rect 0 37408 800 37528
rect 179200 33192 180000 33312
rect 0 32376 800 32496
rect 179200 28840 180000 28960
rect 0 27344 800 27464
rect 179200 24352 180000 24472
rect 0 22448 800 22568
rect 179200 19864 180000 19984
rect 0 17416 800 17536
rect 179200 15512 180000 15632
rect 0 12384 800 12504
rect 179200 11024 180000 11144
rect 0 7352 800 7472
rect 179200 6536 180000 6656
rect 0 2456 800 2576
rect 179200 2184 180000 2304
<< obsm3 >>
rect 880 117296 179200 117537
rect 800 113360 179200 117296
rect 800 113080 179120 113360
rect 800 112544 179200 113080
rect 880 112264 179200 112544
rect 800 109008 179200 112264
rect 800 108728 179120 109008
rect 800 107512 179200 108728
rect 880 107232 179200 107512
rect 800 104520 179200 107232
rect 800 104240 179120 104520
rect 800 102616 179200 104240
rect 880 102336 179200 102616
rect 800 100032 179200 102336
rect 800 99752 179120 100032
rect 800 97584 179200 99752
rect 880 97304 179200 97584
rect 800 95680 179200 97304
rect 800 95400 179120 95680
rect 800 92552 179200 95400
rect 880 92272 179200 92552
rect 800 91192 179200 92272
rect 800 90912 179120 91192
rect 800 87520 179200 90912
rect 880 87240 179200 87520
rect 800 86704 179200 87240
rect 800 86424 179120 86704
rect 800 82624 179200 86424
rect 880 82352 179200 82624
rect 880 82344 179120 82352
rect 800 82072 179120 82344
rect 800 77864 179200 82072
rect 800 77592 179120 77864
rect 880 77584 179120 77592
rect 880 77312 179200 77584
rect 800 73376 179200 77312
rect 800 73096 179120 73376
rect 800 72560 179200 73096
rect 880 72280 179200 72560
rect 800 69024 179200 72280
rect 800 68744 179120 69024
rect 800 67528 179200 68744
rect 880 67248 179200 67528
rect 800 64536 179200 67248
rect 800 64256 179120 64536
rect 800 62632 179200 64256
rect 880 62352 179200 62632
rect 800 60048 179200 62352
rect 800 59768 179120 60048
rect 800 57600 179200 59768
rect 880 57320 179200 57600
rect 800 55696 179200 57320
rect 800 55416 179120 55696
rect 800 52568 179200 55416
rect 880 52288 179200 52568
rect 800 51208 179200 52288
rect 800 50928 179120 51208
rect 800 47536 179200 50928
rect 880 47256 179200 47536
rect 800 46720 179200 47256
rect 800 46440 179120 46720
rect 800 42640 179200 46440
rect 880 42368 179200 42640
rect 880 42360 179120 42368
rect 800 42088 179120 42360
rect 800 37880 179200 42088
rect 800 37608 179120 37880
rect 880 37600 179120 37608
rect 880 37328 179200 37600
rect 800 33392 179200 37328
rect 800 33112 179120 33392
rect 800 32576 179200 33112
rect 880 32296 179200 32576
rect 800 29040 179200 32296
rect 800 28760 179120 29040
rect 800 27544 179200 28760
rect 880 27264 179200 27544
rect 800 24552 179200 27264
rect 800 24272 179120 24552
rect 800 22648 179200 24272
rect 880 22368 179200 22648
rect 800 20064 179200 22368
rect 800 19784 179120 20064
rect 800 17616 179200 19784
rect 880 17336 179200 17616
rect 800 15712 179200 17336
rect 800 15432 179120 15712
rect 800 12584 179200 15432
rect 880 12304 179200 12584
rect 800 11224 179200 12304
rect 800 10944 179120 11224
rect 800 7552 179200 10944
rect 880 7272 179200 7552
rect 800 6736 179200 7272
rect 800 6456 179120 6736
rect 800 2656 179200 6456
rect 880 2384 179200 2656
rect 880 2376 179120 2384
rect 800 2143 179120 2376
<< metal4 >>
rect 4208 2128 4528 117552
rect 19568 2128 19888 117552
rect 34928 2128 35248 117552
rect 50288 2128 50608 117552
rect 65648 2128 65968 117552
rect 81008 2128 81328 117552
rect 96368 2128 96688 117552
rect 111728 2128 112048 117552
rect 127088 2128 127408 117552
rect 142448 2128 142768 117552
rect 157808 2128 158128 117552
rect 173168 2128 173488 117552
<< obsm4 >>
rect 99051 114411 99117 117333
<< labels >>
rlabel metal2 s 33690 0 33746 800 6 addr0[0]
port 1 nsew signal input
rlabel metal3 s 179200 68824 180000 68944 6 addr0[10]
port 2 nsew signal input
rlabel metal3 s 179200 77664 180000 77784 6 addr0[11]
port 3 nsew signal input
rlabel metal3 s 179200 86504 180000 86624 6 addr0[12]
port 4 nsew signal input
rlabel metal3 s 0 77392 800 77512 6 addr0[13]
port 5 nsew signal input
rlabel metal2 s 153934 119200 153990 120000 6 addr0[14]
port 6 nsew signal input
rlabel metal3 s 0 97384 800 97504 6 addr0[15]
port 7 nsew signal input
rlabel metal3 s 0 107312 800 107432 6 addr0[16]
port 8 nsew signal input
rlabel metal3 s 0 112344 800 112464 6 addr0[17]
port 9 nsew signal input
rlabel metal3 s 179200 95480 180000 95600 6 addr0[18]
port 10 nsew signal input
rlabel metal2 s 158626 119200 158682 120000 6 addr0[19]
port 11 nsew signal input
rlabel metal3 s 0 12384 800 12504 6 addr0[1]
port 12 nsew signal input
rlabel metal2 s 168654 0 168710 800 6 addr0[20]
port 13 nsew signal input
rlabel metal2 s 163410 119200 163466 120000 6 addr0[21]
port 14 nsew signal input
rlabel metal2 s 168102 119200 168158 120000 6 addr0[22]
port 15 nsew signal input
rlabel metal3 s 179200 99832 180000 99952 6 addr0[23]
port 16 nsew signal input
rlabel metal3 s 0 117376 800 117496 6 addr0[24]
port 17 nsew signal input
rlabel metal2 s 176198 0 176254 800 6 addr0[25]
port 18 nsew signal input
rlabel metal3 s 179200 104320 180000 104440 6 addr0[26]
port 19 nsew signal input
rlabel metal2 s 172886 119200 172942 120000 6 addr0[27]
port 20 nsew signal input
rlabel metal3 s 179200 108808 180000 108928 6 addr0[28]
port 21 nsew signal input
rlabel metal3 s 179200 113160 180000 113280 6 addr0[29]
port 22 nsew signal input
rlabel metal2 s 78678 0 78734 800 6 addr0[2]
port 23 nsew signal input
rlabel metal2 s 177578 119200 177634 120000 6 addr0[30]
port 24 nsew signal input
rlabel metal3 s 179200 117648 180000 117768 6 addr0[31]
port 25 nsew signal input
rlabel metal3 s 0 22448 800 22568 6 addr0[3]
port 26 nsew signal input
rlabel metal3 s 0 27344 800 27464 6 addr0[4]
port 27 nsew signal input
rlabel metal3 s 0 47336 800 47456 6 addr0[5]
port 28 nsew signal input
rlabel metal2 s 116214 0 116270 800 6 addr0[6]
port 29 nsew signal input
rlabel metal3 s 179200 46520 180000 46640 6 addr0[7]
port 30 nsew signal input
rlabel metal3 s 179200 55496 180000 55616 6 addr0[8]
port 31 nsew signal input
rlabel metal3 s 179200 64336 180000 64456 6 addr0[9]
port 32 nsew signal input
rlabel metal3 s 0 2456 800 2576 6 b
port 33 nsew signal output
rlabel metal2 s 101770 119200 101826 120000 6 clk
port 34 nsew signal input
rlabel metal3 s 179200 2184 180000 2304 6 din0[0]
port 35 nsew signal input
rlabel metal2 s 146206 0 146262 800 6 din0[10]
port 36 nsew signal input
rlabel metal3 s 179200 82152 180000 82272 6 din0[11]
port 37 nsew signal input
rlabel metal2 s 149150 119200 149206 120000 6 din0[12]
port 38 nsew signal input
rlabel metal3 s 0 82424 800 82544 6 din0[13]
port 39 nsew signal input
rlabel metal3 s 0 92352 800 92472 6 din0[14]
port 40 nsew signal input
rlabel metal3 s 0 102416 800 102536 6 din0[15]
port 41 nsew signal input
rlabel metal3 s 0 17416 800 17536 6 din0[1]
port 42 nsew signal input
rlabel metal2 s 134982 119200 135038 120000 6 din0[2]
port 43 nsew signal input
rlabel metal3 s 179200 15512 180000 15632 6 din0[3]
port 44 nsew signal input
rlabel metal3 s 0 32376 800 32496 6 din0[4]
port 45 nsew signal input
rlabel metal2 s 101218 0 101274 800 6 din0[5]
port 46 nsew signal input
rlabel metal2 s 123666 0 123722 800 6 din0[6]
port 47 nsew signal input
rlabel metal3 s 0 57400 800 57520 6 din0[7]
port 48 nsew signal input
rlabel metal3 s 179200 59848 180000 59968 6 din0[8]
port 49 nsew signal input
rlabel metal3 s 0 67328 800 67448 6 din0[9]
port 50 nsew signal input
rlabel metal3 s 0 7352 800 7472 6 din[0]
port 51 nsew signal input
rlabel metal2 s 56138 0 56194 800 6 din[1]
port 52 nsew signal input
rlabel metal2 s 86130 0 86186 800 6 din[2]
port 53 nsew signal input
rlabel metal3 s 179200 19864 180000 19984 6 din[3]
port 54 nsew signal input
rlabel metal3 s 0 37408 800 37528 6 din[4]
port 55 nsew signal input
rlabel metal3 s 179200 28840 180000 28960 6 din[5]
port 56 nsew signal input
rlabel metal3 s 179200 37680 180000 37800 6 din[6]
port 57 nsew signal input
rlabel metal3 s 179200 51008 180000 51128 6 din[7]
port 58 nsew signal input
rlabel metal2 s 41142 0 41198 800 6 dout0[0]
port 59 nsew signal output
rlabel metal3 s 179200 73176 180000 73296 6 dout0[10]
port 60 nsew signal output
rlabel metal3 s 0 72360 800 72480 6 dout0[11]
port 61 nsew signal output
rlabel metal3 s 179200 90992 180000 91112 6 dout0[12]
port 62 nsew signal output
rlabel metal3 s 0 87320 800 87440 6 dout0[13]
port 63 nsew signal output
rlabel metal2 s 153658 0 153714 800 6 dout0[14]
port 64 nsew signal output
rlabel metal2 s 161202 0 161258 800 6 dout0[15]
port 65 nsew signal output
rlabel metal2 s 63682 0 63738 800 6 dout0[1]
port 66 nsew signal output
rlabel metal3 s 179200 6536 180000 6656 6 dout0[2]
port 67 nsew signal output
rlabel metal3 s 179200 24352 180000 24472 6 dout0[3]
port 68 nsew signal output
rlabel metal2 s 93674 0 93730 800 6 dout0[4]
port 69 nsew signal output
rlabel metal3 s 179200 33192 180000 33312 6 dout0[5]
port 70 nsew signal output
rlabel metal3 s 0 52368 800 52488 6 dout0[6]
port 71 nsew signal output
rlabel metal3 s 0 62432 800 62552 6 dout0[7]
port 72 nsew signal output
rlabel metal2 s 144458 119200 144514 120000 6 dout0[8]
port 73 nsew signal output
rlabel metal2 s 138662 0 138718 800 6 dout0[9]
port 74 nsew signal output
rlabel metal2 s 48686 0 48742 800 6 dout[0]
port 75 nsew signal output
rlabel metal2 s 130198 119200 130254 120000 6 dout[1]
port 76 nsew signal output
rlabel metal3 s 179200 11024 180000 11144 6 dout[2]
port 77 nsew signal output
rlabel metal2 s 139674 119200 139730 120000 6 dout[3]
port 78 nsew signal output
rlabel metal3 s 0 42440 800 42560 6 dout[4]
port 79 nsew signal output
rlabel metal2 s 108670 0 108726 800 6 dout[5]
port 80 nsew signal output
rlabel metal3 s 179200 42168 180000 42288 6 dout[6]
port 81 nsew signal output
rlabel metal2 s 131210 0 131266 800 6 dout[7]
port 82 nsew signal output
rlabel metal2 s 18694 0 18750 800 6 g
port 83 nsew signal output
rlabel metal2 s 106554 119200 106610 120000 6 hs
port 84 nsew signal output
rlabel metal2 s 2318 119200 2374 120000 6 io_oeb[0]
port 85 nsew signal output
rlabel metal2 s 49698 119200 49754 120000 6 io_oeb[10]
port 86 nsew signal output
rlabel metal2 s 54390 119200 54446 120000 6 io_oeb[11]
port 87 nsew signal output
rlabel metal2 s 59174 119200 59230 120000 6 io_oeb[12]
port 88 nsew signal output
rlabel metal2 s 63866 119200 63922 120000 6 io_oeb[13]
port 89 nsew signal output
rlabel metal2 s 68650 119200 68706 120000 6 io_oeb[14]
port 90 nsew signal output
rlabel metal2 s 73342 119200 73398 120000 6 io_oeb[15]
port 91 nsew signal output
rlabel metal2 s 78126 119200 78182 120000 6 io_oeb[16]
port 92 nsew signal output
rlabel metal2 s 82818 119200 82874 120000 6 io_oeb[17]
port 93 nsew signal output
rlabel metal2 s 87602 119200 87658 120000 6 io_oeb[18]
port 94 nsew signal output
rlabel metal2 s 92294 119200 92350 120000 6 io_oeb[19]
port 95 nsew signal output
rlabel metal2 s 7010 119200 7066 120000 6 io_oeb[1]
port 96 nsew signal output
rlabel metal2 s 97078 119200 97134 120000 6 io_oeb[20]
port 97 nsew signal output
rlabel metal2 s 11794 119200 11850 120000 6 io_oeb[2]
port 98 nsew signal output
rlabel metal2 s 16486 119200 16542 120000 6 io_oeb[3]
port 99 nsew signal output
rlabel metal2 s 21270 119200 21326 120000 6 io_oeb[4]
port 100 nsew signal output
rlabel metal2 s 25962 119200 26018 120000 6 io_oeb[5]
port 101 nsew signal output
rlabel metal2 s 30746 119200 30802 120000 6 io_oeb[6]
port 102 nsew signal output
rlabel metal2 s 35438 119200 35494 120000 6 io_oeb[7]
port 103 nsew signal output
rlabel metal2 s 40222 119200 40278 120000 6 io_oeb[8]
port 104 nsew signal output
rlabel metal2 s 44914 119200 44970 120000 6 io_oeb[9]
port 105 nsew signal output
rlabel metal2 s 26146 0 26202 800 6 r
port 106 nsew signal output
rlabel metal2 s 111246 119200 111302 120000 6 rst
port 107 nsew signal input
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 108 nsew power input
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 108 nsew power input
rlabel metal4 s 65648 2128 65968 117552 6 vccd1
port 108 nsew power input
rlabel metal4 s 96368 2128 96688 117552 6 vccd1
port 108 nsew power input
rlabel metal4 s 127088 2128 127408 117552 6 vccd1
port 108 nsew power input
rlabel metal4 s 157808 2128 158128 117552 6 vccd1
port 108 nsew power input
rlabel metal2 s 116030 119200 116086 120000 6 vs
port 109 nsew signal output
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 110 nsew ground input
rlabel metal4 s 50288 2128 50608 117552 6 vssd1
port 110 nsew ground input
rlabel metal4 s 81008 2128 81328 117552 6 vssd1
port 110 nsew ground input
rlabel metal4 s 111728 2128 112048 117552 6 vssd1
port 110 nsew ground input
rlabel metal4 s 142448 2128 142768 117552 6 vssd1
port 110 nsew ground input
rlabel metal4 s 173168 2128 173488 117552 6 vssd1
port 110 nsew ground input
rlabel metal2 s 3698 0 3754 800 6 wbs_cyc_i
port 111 nsew signal input
rlabel metal2 s 11150 0 11206 800 6 wbs_stb_i
port 112 nsew signal input
rlabel metal2 s 120722 119200 120778 120000 6 web
port 113 nsew signal input
rlabel metal2 s 125506 119200 125562 120000 6 wmask0[0]
port 114 nsew signal input
rlabel metal2 s 71134 0 71190 800 6 wmask0[1]
port 115 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 180000 120000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 6006776
string GDS_FILE /home/fabio/chip_tutorial/upb_natalius_soc/openlane/natalius_soc/runs/natalius_soc/results/finishing/natalius_soc.magic.gds
string GDS_START 263090
<< end >>

