VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO natalius_soc
  CLASS BLOCK ;
  FOREIGN natalius_soc ;
  ORIGIN 0.000 0.000 ;
  SIZE 900.000 BY 600.000 ;
  PIN addr0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.450 0.000 168.730 4.000 ;
    END
  END addr0[0]
  PIN addr0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 344.120 900.000 344.720 ;
    END
  END addr0[10]
  PIN addr0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 388.320 900.000 388.920 ;
    END
  END addr0[11]
  PIN addr0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 432.520 900.000 433.120 ;
    END
  END addr0[12]
  PIN addr0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 386.960 4.000 387.560 ;
    END
  END addr0[13]
  PIN addr0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 769.670 596.000 769.950 600.000 ;
    END
  END addr0[14]
  PIN addr0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 486.920 4.000 487.520 ;
    END
  END addr0[15]
  PIN addr0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 536.560 4.000 537.160 ;
    END
  END addr0[16]
  PIN addr0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 561.720 4.000 562.320 ;
    END
  END addr0[17]
  PIN addr0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 477.400 900.000 478.000 ;
    END
  END addr0[18]
  PIN addr0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 793.130 596.000 793.410 600.000 ;
    END
  END addr0[19]
  PIN addr0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.920 4.000 62.520 ;
    END
  END addr0[1]
  PIN addr0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 843.270 0.000 843.550 4.000 ;
    END
  END addr0[20]
  PIN addr0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 817.050 596.000 817.330 600.000 ;
    END
  END addr0[21]
  PIN addr0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 840.510 596.000 840.790 600.000 ;
    END
  END addr0[22]
  PIN addr0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 499.160 900.000 499.760 ;
    END
  END addr0[23]
  PIN addr0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 586.880 4.000 587.480 ;
    END
  END addr0[24]
  PIN addr0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 880.990 0.000 881.270 4.000 ;
    END
  END addr0[25]
  PIN addr0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 521.600 900.000 522.200 ;
    END
  END addr0[26]
  PIN addr0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 864.430 596.000 864.710 600.000 ;
    END
  END addr0[27]
  PIN addr0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 544.040 900.000 544.640 ;
    END
  END addr0[28]
  PIN addr0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 565.800 900.000 566.400 ;
    END
  END addr0[29]
  PIN addr0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.390 0.000 393.670 4.000 ;
    END
  END addr0[2]
  PIN addr0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 887.890 596.000 888.170 600.000 ;
    END
  END addr0[30]
  PIN addr0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 588.240 900.000 588.840 ;
    END
  END addr0[31]
  PIN addr0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 4.000 112.840 ;
    END
  END addr0[3]
  PIN addr0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.720 4.000 137.320 ;
    END
  END addr0[4]
  PIN addr0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 236.680 4.000 237.280 ;
    END
  END addr0[5]
  PIN addr0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.070 0.000 581.350 4.000 ;
    END
  END addr0[6]
  PIN addr0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 232.600 900.000 233.200 ;
    END
  END addr0[7]
  PIN addr0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 277.480 900.000 278.080 ;
    END
  END addr0[8]
  PIN addr0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 321.680 900.000 322.280 ;
    END
  END addr0[9]
  PIN b
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.280 4.000 12.880 ;
    END
  END b
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.850 596.000 509.130 600.000 ;
    END
  END clk
  PIN din0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 10.920 900.000 11.520 ;
    END
  END din0[0]
  PIN din0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 731.030 0.000 731.310 4.000 ;
    END
  END din0[10]
  PIN din0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 410.760 900.000 411.360 ;
    END
  END din0[11]
  PIN din0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 745.750 596.000 746.030 600.000 ;
    END
  END din0[12]
  PIN din0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 412.120 4.000 412.720 ;
    END
  END din0[13]
  PIN din0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 461.760 4.000 462.360 ;
    END
  END din0[14]
  PIN din0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 512.080 4.000 512.680 ;
    END
  END din0[15]
  PIN din0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.080 4.000 87.680 ;
    END
  END din0[1]
  PIN din0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 674.910 596.000 675.190 600.000 ;
    END
  END din0[2]
  PIN din0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 77.560 900.000 78.160 ;
    END
  END din0[3]
  PIN din0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.880 4.000 162.480 ;
    END
  END din0[4]
  PIN din0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 506.090 0.000 506.370 4.000 ;
    END
  END din0[5]
  PIN din0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 618.330 0.000 618.610 4.000 ;
    END
  END din0[6]
  PIN din0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 287.000 4.000 287.600 ;
    END
  END din0[7]
  PIN din0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 299.240 900.000 299.840 ;
    END
  END din0[8]
  PIN din0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 336.640 4.000 337.240 ;
    END
  END din0[9]
  PIN din[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.760 4.000 37.360 ;
    END
  END din[0]
  PIN din[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.690 0.000 280.970 4.000 ;
    END
  END din[1]
  PIN din[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.650 0.000 430.930 4.000 ;
    END
  END din[2]
  PIN din[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 99.320 900.000 99.920 ;
    END
  END din[3]
  PIN din[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.040 4.000 187.640 ;
    END
  END din[4]
  PIN din[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 144.200 900.000 144.800 ;
    END
  END din[5]
  PIN din[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 188.400 900.000 189.000 ;
    END
  END din[6]
  PIN din[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 255.040 900.000 255.640 ;
    END
  END din[7]
  PIN dout0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.710 0.000 205.990 4.000 ;
    END
  END dout0[0]
  PIN dout0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 365.880 900.000 366.480 ;
    END
  END dout0[10]
  PIN dout0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 361.800 4.000 362.400 ;
    END
  END dout0[11]
  PIN dout0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 454.960 900.000 455.560 ;
    END
  END dout0[12]
  PIN dout0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 436.600 4.000 437.200 ;
    END
  END dout0[13]
  PIN dout0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 768.290 0.000 768.570 4.000 ;
    END
  END dout0[14]
  PIN dout0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 806.010 0.000 806.290 4.000 ;
    END
  END dout0[15]
  PIN dout0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.410 0.000 318.690 4.000 ;
    END
  END dout0[1]
  PIN dout0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 32.680 900.000 33.280 ;
    END
  END dout0[2]
  PIN dout0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 121.760 900.000 122.360 ;
    END
  END dout0[3]
  PIN dout0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 468.370 0.000 468.650 4.000 ;
    END
  END dout0[4]
  PIN dout0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 165.960 900.000 166.560 ;
    END
  END dout0[5]
  PIN dout0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.840 4.000 262.440 ;
    END
  END dout0[6]
  PIN dout0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.160 4.000 312.760 ;
    END
  END dout0[7]
  PIN dout0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 722.290 596.000 722.570 600.000 ;
    END
  END dout0[8]
  PIN dout0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 693.310 0.000 693.590 4.000 ;
    END
  END dout0[9]
  PIN dout[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.430 0.000 243.710 4.000 ;
    END
  END dout[0]
  PIN dout[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.990 596.000 651.270 600.000 ;
    END
  END dout[1]
  PIN dout[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 55.120 900.000 55.720 ;
    END
  END dout[2]
  PIN dout[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 698.370 596.000 698.650 600.000 ;
    END
  END dout[3]
  PIN dout[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.200 4.000 212.800 ;
    END
  END dout[4]
  PIN dout[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 543.350 0.000 543.630 4.000 ;
    END
  END dout[5]
  PIN dout[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 210.840 900.000 211.440 ;
    END
  END dout[6]
  PIN dout[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.050 0.000 656.330 4.000 ;
    END
  END dout[7]
  PIN g
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 4.000 ;
    END
  END g
  PIN hs
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 532.770 596.000 533.050 600.000 ;
    END
  END hs
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 596.000 11.870 600.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.490 596.000 248.770 600.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.950 596.000 272.230 600.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 295.870 596.000 296.150 600.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.330 596.000 319.610 600.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.250 596.000 343.530 600.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.710 596.000 366.990 600.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.630 596.000 390.910 600.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.090 596.000 414.370 600.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.010 596.000 438.290 600.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.470 596.000 461.750 600.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.050 596.000 35.330 600.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 485.390 596.000 485.670 600.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.970 596.000 59.250 600.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.430 596.000 82.710 600.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 596.000 106.630 600.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.810 596.000 130.090 600.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.730 596.000 154.010 600.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 596.000 177.470 600.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.110 596.000 201.390 600.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.570 596.000 224.850 600.000 ;
    END
  END io_oeb[9]
  PIN r
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.730 0.000 131.010 4.000 ;
    END
  END r
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.230 596.000 556.510 600.000 ;
    END
  END rst
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 587.760 ;
    END
  END vccd1
  PIN vs
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 580.150 596.000 580.430 600.000 ;
    END
  END vs
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 587.760 ;
    END
  END vssd1
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.490 0.000 18.770 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 0.000 56.030 4.000 ;
    END
  END wbs_stb_i
  PIN web
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 603.610 596.000 603.890 600.000 ;
    END
  END web
  PIN wmask0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.530 596.000 627.810 600.000 ;
    END
  END wmask0[0]
  PIN wmask0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 355.670 0.000 355.950 4.000 ;
    END
  END wmask0[1]
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 894.240 587.605 ;
      LAYER met1 ;
        RECT 5.520 10.640 894.240 589.520 ;
      LAYER met2 ;
        RECT 6.990 595.720 11.310 596.770 ;
        RECT 12.150 595.720 34.770 596.770 ;
        RECT 35.610 595.720 58.690 596.770 ;
        RECT 59.530 595.720 82.150 596.770 ;
        RECT 82.990 595.720 106.070 596.770 ;
        RECT 106.910 595.720 129.530 596.770 ;
        RECT 130.370 595.720 153.450 596.770 ;
        RECT 154.290 595.720 176.910 596.770 ;
        RECT 177.750 595.720 200.830 596.770 ;
        RECT 201.670 595.720 224.290 596.770 ;
        RECT 225.130 595.720 248.210 596.770 ;
        RECT 249.050 595.720 271.670 596.770 ;
        RECT 272.510 595.720 295.590 596.770 ;
        RECT 296.430 595.720 319.050 596.770 ;
        RECT 319.890 595.720 342.970 596.770 ;
        RECT 343.810 595.720 366.430 596.770 ;
        RECT 367.270 595.720 390.350 596.770 ;
        RECT 391.190 595.720 413.810 596.770 ;
        RECT 414.650 595.720 437.730 596.770 ;
        RECT 438.570 595.720 461.190 596.770 ;
        RECT 462.030 595.720 485.110 596.770 ;
        RECT 485.950 595.720 508.570 596.770 ;
        RECT 509.410 595.720 532.490 596.770 ;
        RECT 533.330 595.720 555.950 596.770 ;
        RECT 556.790 595.720 579.870 596.770 ;
        RECT 580.710 595.720 603.330 596.770 ;
        RECT 604.170 595.720 627.250 596.770 ;
        RECT 628.090 595.720 650.710 596.770 ;
        RECT 651.550 595.720 674.630 596.770 ;
        RECT 675.470 595.720 698.090 596.770 ;
        RECT 698.930 595.720 722.010 596.770 ;
        RECT 722.850 595.720 745.470 596.770 ;
        RECT 746.310 595.720 769.390 596.770 ;
        RECT 770.230 595.720 792.850 596.770 ;
        RECT 793.690 595.720 816.770 596.770 ;
        RECT 817.610 595.720 840.230 596.770 ;
        RECT 841.070 595.720 864.150 596.770 ;
        RECT 864.990 595.720 887.610 596.770 ;
        RECT 888.450 595.720 890.930 596.770 ;
        RECT 6.990 4.280 890.930 595.720 ;
        RECT 6.990 4.000 18.210 4.280 ;
        RECT 19.050 4.000 55.470 4.280 ;
        RECT 56.310 4.000 93.190 4.280 ;
        RECT 94.030 4.000 130.450 4.280 ;
        RECT 131.290 4.000 168.170 4.280 ;
        RECT 169.010 4.000 205.430 4.280 ;
        RECT 206.270 4.000 243.150 4.280 ;
        RECT 243.990 4.000 280.410 4.280 ;
        RECT 281.250 4.000 318.130 4.280 ;
        RECT 318.970 4.000 355.390 4.280 ;
        RECT 356.230 4.000 393.110 4.280 ;
        RECT 393.950 4.000 430.370 4.280 ;
        RECT 431.210 4.000 468.090 4.280 ;
        RECT 468.930 4.000 505.810 4.280 ;
        RECT 506.650 4.000 543.070 4.280 ;
        RECT 543.910 4.000 580.790 4.280 ;
        RECT 581.630 4.000 618.050 4.280 ;
        RECT 618.890 4.000 655.770 4.280 ;
        RECT 656.610 4.000 693.030 4.280 ;
        RECT 693.870 4.000 730.750 4.280 ;
        RECT 731.590 4.000 768.010 4.280 ;
        RECT 768.850 4.000 805.730 4.280 ;
        RECT 806.570 4.000 842.990 4.280 ;
        RECT 843.830 4.000 880.710 4.280 ;
        RECT 881.550 4.000 890.930 4.280 ;
      LAYER met3 ;
        RECT 4.400 586.480 896.000 587.685 ;
        RECT 4.000 566.800 896.000 586.480 ;
        RECT 4.000 565.400 895.600 566.800 ;
        RECT 4.000 562.720 896.000 565.400 ;
        RECT 4.400 561.320 896.000 562.720 ;
        RECT 4.000 545.040 896.000 561.320 ;
        RECT 4.000 543.640 895.600 545.040 ;
        RECT 4.000 537.560 896.000 543.640 ;
        RECT 4.400 536.160 896.000 537.560 ;
        RECT 4.000 522.600 896.000 536.160 ;
        RECT 4.000 521.200 895.600 522.600 ;
        RECT 4.000 513.080 896.000 521.200 ;
        RECT 4.400 511.680 896.000 513.080 ;
        RECT 4.000 500.160 896.000 511.680 ;
        RECT 4.000 498.760 895.600 500.160 ;
        RECT 4.000 487.920 896.000 498.760 ;
        RECT 4.400 486.520 896.000 487.920 ;
        RECT 4.000 478.400 896.000 486.520 ;
        RECT 4.000 477.000 895.600 478.400 ;
        RECT 4.000 462.760 896.000 477.000 ;
        RECT 4.400 461.360 896.000 462.760 ;
        RECT 4.000 455.960 896.000 461.360 ;
        RECT 4.000 454.560 895.600 455.960 ;
        RECT 4.000 437.600 896.000 454.560 ;
        RECT 4.400 436.200 896.000 437.600 ;
        RECT 4.000 433.520 896.000 436.200 ;
        RECT 4.000 432.120 895.600 433.520 ;
        RECT 4.000 413.120 896.000 432.120 ;
        RECT 4.400 411.760 896.000 413.120 ;
        RECT 4.400 411.720 895.600 411.760 ;
        RECT 4.000 410.360 895.600 411.720 ;
        RECT 4.000 389.320 896.000 410.360 ;
        RECT 4.000 387.960 895.600 389.320 ;
        RECT 4.400 387.920 895.600 387.960 ;
        RECT 4.400 386.560 896.000 387.920 ;
        RECT 4.000 366.880 896.000 386.560 ;
        RECT 4.000 365.480 895.600 366.880 ;
        RECT 4.000 362.800 896.000 365.480 ;
        RECT 4.400 361.400 896.000 362.800 ;
        RECT 4.000 345.120 896.000 361.400 ;
        RECT 4.000 343.720 895.600 345.120 ;
        RECT 4.000 337.640 896.000 343.720 ;
        RECT 4.400 336.240 896.000 337.640 ;
        RECT 4.000 322.680 896.000 336.240 ;
        RECT 4.000 321.280 895.600 322.680 ;
        RECT 4.000 313.160 896.000 321.280 ;
        RECT 4.400 311.760 896.000 313.160 ;
        RECT 4.000 300.240 896.000 311.760 ;
        RECT 4.000 298.840 895.600 300.240 ;
        RECT 4.000 288.000 896.000 298.840 ;
        RECT 4.400 286.600 896.000 288.000 ;
        RECT 4.000 278.480 896.000 286.600 ;
        RECT 4.000 277.080 895.600 278.480 ;
        RECT 4.000 262.840 896.000 277.080 ;
        RECT 4.400 261.440 896.000 262.840 ;
        RECT 4.000 256.040 896.000 261.440 ;
        RECT 4.000 254.640 895.600 256.040 ;
        RECT 4.000 237.680 896.000 254.640 ;
        RECT 4.400 236.280 896.000 237.680 ;
        RECT 4.000 233.600 896.000 236.280 ;
        RECT 4.000 232.200 895.600 233.600 ;
        RECT 4.000 213.200 896.000 232.200 ;
        RECT 4.400 211.840 896.000 213.200 ;
        RECT 4.400 211.800 895.600 211.840 ;
        RECT 4.000 210.440 895.600 211.800 ;
        RECT 4.000 189.400 896.000 210.440 ;
        RECT 4.000 188.040 895.600 189.400 ;
        RECT 4.400 188.000 895.600 188.040 ;
        RECT 4.400 186.640 896.000 188.000 ;
        RECT 4.000 166.960 896.000 186.640 ;
        RECT 4.000 165.560 895.600 166.960 ;
        RECT 4.000 162.880 896.000 165.560 ;
        RECT 4.400 161.480 896.000 162.880 ;
        RECT 4.000 145.200 896.000 161.480 ;
        RECT 4.000 143.800 895.600 145.200 ;
        RECT 4.000 137.720 896.000 143.800 ;
        RECT 4.400 136.320 896.000 137.720 ;
        RECT 4.000 122.760 896.000 136.320 ;
        RECT 4.000 121.360 895.600 122.760 ;
        RECT 4.000 113.240 896.000 121.360 ;
        RECT 4.400 111.840 896.000 113.240 ;
        RECT 4.000 100.320 896.000 111.840 ;
        RECT 4.000 98.920 895.600 100.320 ;
        RECT 4.000 88.080 896.000 98.920 ;
        RECT 4.400 86.680 896.000 88.080 ;
        RECT 4.000 78.560 896.000 86.680 ;
        RECT 4.000 77.160 895.600 78.560 ;
        RECT 4.000 62.920 896.000 77.160 ;
        RECT 4.400 61.520 896.000 62.920 ;
        RECT 4.000 56.120 896.000 61.520 ;
        RECT 4.000 54.720 895.600 56.120 ;
        RECT 4.000 37.760 896.000 54.720 ;
        RECT 4.400 36.360 896.000 37.760 ;
        RECT 4.000 33.680 896.000 36.360 ;
        RECT 4.000 32.280 895.600 33.680 ;
        RECT 4.000 13.280 896.000 32.280 ;
        RECT 4.400 11.920 896.000 13.280 ;
        RECT 4.400 11.880 895.600 11.920 ;
        RECT 4.000 10.715 895.600 11.880 ;
      LAYER met4 ;
        RECT 495.255 572.055 495.585 586.665 ;
  END
END natalius_soc
END LIBRARY

