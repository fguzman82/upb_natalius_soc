magic
tech sky130A
magscale 1 2
timestamp 1654745837
<< obsli1 >>
rect 1104 2159 178848 117521
<< obsm1 >>
rect 1104 2128 178848 117552
<< metal2 >>
rect 2134 119200 2190 120000
rect 6366 119200 6422 120000
rect 10690 119200 10746 120000
rect 14922 119200 14978 120000
rect 19246 119200 19302 120000
rect 23478 119200 23534 120000
rect 27802 119200 27858 120000
rect 32126 119200 32182 120000
rect 36358 119200 36414 120000
rect 40682 119200 40738 120000
rect 44914 119200 44970 120000
rect 49238 119200 49294 120000
rect 53562 119200 53618 120000
rect 57794 119200 57850 120000
rect 62118 119200 62174 120000
rect 66350 119200 66406 120000
rect 70674 119200 70730 120000
rect 74998 119200 75054 120000
rect 79230 119200 79286 120000
rect 83554 119200 83610 120000
rect 87786 119200 87842 120000
rect 92110 119200 92166 120000
rect 96434 119200 96490 120000
rect 100666 119200 100722 120000
rect 104990 119200 105046 120000
rect 109222 119200 109278 120000
rect 113546 119200 113602 120000
rect 117870 119200 117926 120000
rect 122102 119200 122158 120000
rect 126426 119200 126482 120000
rect 130658 119200 130714 120000
rect 134982 119200 135038 120000
rect 139306 119200 139362 120000
rect 143538 119200 143594 120000
rect 147862 119200 147918 120000
rect 152094 119200 152150 120000
rect 156418 119200 156474 120000
rect 160742 119200 160798 120000
rect 164974 119200 165030 120000
rect 169298 119200 169354 120000
rect 173530 119200 173586 120000
rect 177854 119200 177910 120000
rect 4066 0 4122 800
rect 12162 0 12218 800
rect 20350 0 20406 800
rect 28538 0 28594 800
rect 36726 0 36782 800
rect 44914 0 44970 800
rect 53102 0 53158 800
rect 61290 0 61346 800
rect 69478 0 69534 800
rect 77666 0 77722 800
rect 85854 0 85910 800
rect 94042 0 94098 800
rect 102230 0 102286 800
rect 110418 0 110474 800
rect 118606 0 118662 800
rect 126794 0 126850 800
rect 134982 0 135038 800
rect 143170 0 143226 800
rect 151358 0 151414 800
rect 159546 0 159602 800
rect 167734 0 167790 800
rect 175922 0 175978 800
<< obsm2 >>
rect 1398 119144 2078 119354
rect 2246 119144 6310 119354
rect 6478 119144 10634 119354
rect 10802 119144 14866 119354
rect 15034 119144 19190 119354
rect 19358 119144 23422 119354
rect 23590 119144 27746 119354
rect 27914 119144 32070 119354
rect 32238 119144 36302 119354
rect 36470 119144 40626 119354
rect 40794 119144 44858 119354
rect 45026 119144 49182 119354
rect 49350 119144 53506 119354
rect 53674 119144 57738 119354
rect 57906 119144 62062 119354
rect 62230 119144 66294 119354
rect 66462 119144 70618 119354
rect 70786 119144 74942 119354
rect 75110 119144 79174 119354
rect 79342 119144 83498 119354
rect 83666 119144 87730 119354
rect 87898 119144 92054 119354
rect 92222 119144 96378 119354
rect 96546 119144 100610 119354
rect 100778 119144 104934 119354
rect 105102 119144 109166 119354
rect 109334 119144 113490 119354
rect 113658 119144 117814 119354
rect 117982 119144 122046 119354
rect 122214 119144 126370 119354
rect 126538 119144 130602 119354
rect 130770 119144 134926 119354
rect 135094 119144 139250 119354
rect 139418 119144 143482 119354
rect 143650 119144 147806 119354
rect 147974 119144 152038 119354
rect 152206 119144 156362 119354
rect 156530 119144 160686 119354
rect 160854 119144 164918 119354
rect 165086 119144 169242 119354
rect 169410 119144 173474 119354
rect 173642 119144 177798 119354
rect 177966 119144 178186 119354
rect 1398 856 178186 119144
rect 1398 800 4010 856
rect 4178 800 12106 856
rect 12274 800 20294 856
rect 20462 800 28482 856
rect 28650 800 36670 856
rect 36838 800 44858 856
rect 45026 800 53046 856
rect 53214 800 61234 856
rect 61402 800 69422 856
rect 69590 800 77610 856
rect 77778 800 85798 856
rect 85966 800 93986 856
rect 94154 800 102174 856
rect 102342 800 110362 856
rect 110530 800 118550 856
rect 118718 800 126738 856
rect 126906 800 134926 856
rect 135094 800 143114 856
rect 143282 800 151302 856
rect 151470 800 159490 856
rect 159658 800 167678 856
rect 167846 800 175866 856
rect 176034 800 178186 856
<< metal3 >>
rect 0 116288 800 116408
rect 179200 114792 180000 114912
rect 0 109216 800 109336
rect 179200 104864 180000 104984
rect 0 102144 800 102264
rect 0 95072 800 95192
rect 179200 94800 180000 94920
rect 0 88000 800 88120
rect 179200 84872 180000 84992
rect 0 80928 800 81048
rect 179200 74808 180000 74928
rect 0 73856 800 73976
rect 0 66784 800 66904
rect 179200 64880 180000 65000
rect 0 59848 800 59968
rect 179200 54816 180000 54936
rect 0 52776 800 52896
rect 0 45704 800 45824
rect 179200 44888 180000 45008
rect 0 38632 800 38752
rect 179200 34824 180000 34944
rect 0 31560 800 31680
rect 179200 24896 180000 25016
rect 0 24488 800 24608
rect 0 17416 800 17536
rect 179200 14832 180000 14952
rect 0 10344 800 10464
rect 179200 4904 180000 5024
rect 0 3408 800 3528
<< obsm3 >>
rect 800 116488 179200 117537
rect 880 116208 179200 116488
rect 800 114992 179200 116208
rect 800 114712 179120 114992
rect 800 109416 179200 114712
rect 880 109136 179200 109416
rect 800 105064 179200 109136
rect 800 104784 179120 105064
rect 800 102344 179200 104784
rect 880 102064 179200 102344
rect 800 95272 179200 102064
rect 880 95000 179200 95272
rect 880 94992 179120 95000
rect 800 94720 179120 94992
rect 800 88200 179200 94720
rect 880 87920 179200 88200
rect 800 85072 179200 87920
rect 800 84792 179120 85072
rect 800 81128 179200 84792
rect 880 80848 179200 81128
rect 800 75008 179200 80848
rect 800 74728 179120 75008
rect 800 74056 179200 74728
rect 880 73776 179200 74056
rect 800 66984 179200 73776
rect 880 66704 179200 66984
rect 800 65080 179200 66704
rect 800 64800 179120 65080
rect 800 60048 179200 64800
rect 880 59768 179200 60048
rect 800 55016 179200 59768
rect 800 54736 179120 55016
rect 800 52976 179200 54736
rect 880 52696 179200 52976
rect 800 45904 179200 52696
rect 880 45624 179200 45904
rect 800 45088 179200 45624
rect 800 44808 179120 45088
rect 800 38832 179200 44808
rect 880 38552 179200 38832
rect 800 35024 179200 38552
rect 800 34744 179120 35024
rect 800 31760 179200 34744
rect 880 31480 179200 31760
rect 800 25096 179200 31480
rect 800 24816 179120 25096
rect 800 24688 179200 24816
rect 880 24408 179200 24688
rect 800 17616 179200 24408
rect 880 17336 179200 17616
rect 800 15032 179200 17336
rect 800 14752 179120 15032
rect 800 10544 179200 14752
rect 880 10264 179200 10544
rect 800 5104 179200 10264
rect 800 4824 179120 5104
rect 800 3608 179200 4824
rect 880 3328 179200 3608
rect 800 2143 179200 3328
<< metal4 >>
rect 4208 2128 4528 117552
rect 19568 2128 19888 117552
rect 34928 2128 35248 117552
rect 50288 2128 50608 117552
rect 65648 2128 65968 117552
rect 81008 2128 81328 117552
rect 96368 2128 96688 117552
rect 111728 2128 112048 117552
rect 127088 2128 127408 117552
rect 142448 2128 142768 117552
rect 157808 2128 158128 117552
rect 173168 2128 173488 117552
<< obsm4 >>
rect 13675 13635 19445 21045
<< labels >>
rlabel metal2 s 92110 119200 92166 120000 6 addr0[0]
port 1 nsew signal input
rlabel metal3 s 0 95072 800 95192 6 addr0[10]
port 2 nsew signal input
rlabel metal2 s 167734 0 167790 800 6 addr0[11]
port 3 nsew signal input
rlabel metal3 s 0 38632 800 38752 6 addr0[1]
port 4 nsew signal input
rlabel metal2 s 117870 119200 117926 120000 6 addr0[2]
port 5 nsew signal input
rlabel metal2 s 122102 119200 122158 120000 6 addr0[3]
port 6 nsew signal input
rlabel metal3 s 179200 44888 180000 45008 6 addr0[4]
port 7 nsew signal input
rlabel metal3 s 0 73856 800 73976 6 addr0[5]
port 8 nsew signal input
rlabel metal2 s 134982 119200 135038 120000 6 addr0[6]
port 9 nsew signal input
rlabel metal2 s 126794 0 126850 800 6 addr0[7]
port 10 nsew signal input
rlabel metal2 s 151358 0 151414 800 6 addr0[8]
port 11 nsew signal input
rlabel metal3 s 179200 94800 180000 94920 6 addr0[9]
port 12 nsew signal input
rlabel metal3 s 0 3408 800 3528 6 b
port 13 nsew signal output
rlabel metal3 s 179200 4904 180000 5024 6 clk
port 14 nsew signal input
rlabel metal2 s 28538 0 28594 800 6 din0[0]
port 15 nsew signal input
rlabel metal3 s 0 102144 800 102264 6 din0[10]
port 16 nsew signal input
rlabel metal2 s 156418 119200 156474 120000 6 din0[11]
port 17 nsew signal input
rlabel metal2 s 164974 119200 165030 120000 6 din0[12]
port 18 nsew signal input
rlabel metal3 s 0 116288 800 116408 6 din0[13]
port 19 nsew signal input
rlabel metal2 s 173530 119200 173586 120000 6 din0[14]
port 20 nsew signal input
rlabel metal2 s 177854 119200 177910 120000 6 din0[15]
port 21 nsew signal input
rlabel metal3 s 0 45704 800 45824 6 din0[1]
port 22 nsew signal input
rlabel metal3 s 0 52776 800 52896 6 din0[2]
port 23 nsew signal input
rlabel metal3 s 0 66784 800 66904 6 din0[3]
port 24 nsew signal input
rlabel metal2 s 126426 119200 126482 120000 6 din0[4]
port 25 nsew signal input
rlabel metal3 s 0 80928 800 81048 6 din0[5]
port 26 nsew signal input
rlabel metal2 s 118606 0 118662 800 6 din0[6]
port 27 nsew signal input
rlabel metal2 s 139306 119200 139362 120000 6 din0[7]
port 28 nsew signal input
rlabel metal2 s 143538 119200 143594 120000 6 din0[8]
port 29 nsew signal input
rlabel metal2 s 152094 119200 152150 120000 6 din0[9]
port 30 nsew signal input
rlabel metal2 s 36726 0 36782 800 6 din[0]
port 31 nsew signal input
rlabel metal2 s 104990 119200 105046 120000 6 din[1]
port 32 nsew signal input
rlabel metal3 s 0 59848 800 59968 6 din[2]
port 33 nsew signal input
rlabel metal2 s 61290 0 61346 800 6 din[3]
port 34 nsew signal input
rlabel metal2 s 85854 0 85910 800 6 din[4]
port 35 nsew signal input
rlabel metal2 s 102230 0 102286 800 6 din[5]
port 36 nsew signal input
rlabel metal3 s 179200 64880 180000 65000 6 din[6]
port 37 nsew signal input
rlabel metal3 s 0 88000 800 88120 6 din[7]
port 38 nsew signal input
rlabel metal2 s 96434 119200 96490 120000 6 dout0[0]
port 39 nsew signal output
rlabel metal3 s 0 109216 800 109336 6 dout0[10]
port 40 nsew signal output
rlabel metal2 s 160742 119200 160798 120000 6 dout0[11]
port 41 nsew signal output
rlabel metal2 s 169298 119200 169354 120000 6 dout0[12]
port 42 nsew signal output
rlabel metal2 s 175922 0 175978 800 6 dout0[13]
port 43 nsew signal output
rlabel metal3 s 179200 104864 180000 104984 6 dout0[14]
port 44 nsew signal output
rlabel metal3 s 179200 114792 180000 114912 6 dout0[15]
port 45 nsew signal output
rlabel metal2 s 44914 0 44970 800 6 dout0[1]
port 46 nsew signal output
rlabel metal2 s 53102 0 53158 800 6 dout0[2]
port 47 nsew signal output
rlabel metal2 s 69478 0 69534 800 6 dout0[3]
port 48 nsew signal output
rlabel metal2 s 94042 0 94098 800 6 dout0[4]
port 49 nsew signal output
rlabel metal3 s 179200 54816 180000 54936 6 dout0[5]
port 50 nsew signal output
rlabel metal3 s 179200 74808 180000 74928 6 dout0[6]
port 51 nsew signal output
rlabel metal2 s 134982 0 135038 800 6 dout0[7]
port 52 nsew signal output
rlabel metal2 s 147862 119200 147918 120000 6 dout0[8]
port 53 nsew signal output
rlabel metal2 s 159546 0 159602 800 6 dout0[9]
port 54 nsew signal output
rlabel metal2 s 100666 119200 100722 120000 6 dout[0]
port 55 nsew signal output
rlabel metal2 s 109222 119200 109278 120000 6 dout[1]
port 56 nsew signal output
rlabel metal3 s 179200 34824 180000 34944 6 dout[2]
port 57 nsew signal output
rlabel metal2 s 77666 0 77722 800 6 dout[3]
port 58 nsew signal output
rlabel metal2 s 130658 119200 130714 120000 6 dout[4]
port 59 nsew signal output
rlabel metal2 s 110418 0 110474 800 6 dout[5]
port 60 nsew signal output
rlabel metal3 s 179200 84872 180000 84992 6 dout[6]
port 61 nsew signal output
rlabel metal2 s 143170 0 143226 800 6 dout[7]
port 62 nsew signal output
rlabel metal3 s 0 10344 800 10464 6 g
port 63 nsew signal output
rlabel metal2 s 20350 0 20406 800 6 hs
port 64 nsew signal output
rlabel metal2 s 2134 119200 2190 120000 6 io_oeb[0]
port 65 nsew signal output
rlabel metal2 s 44914 119200 44970 120000 6 io_oeb[10]
port 66 nsew signal output
rlabel metal2 s 49238 119200 49294 120000 6 io_oeb[11]
port 67 nsew signal output
rlabel metal2 s 53562 119200 53618 120000 6 io_oeb[12]
port 68 nsew signal output
rlabel metal2 s 57794 119200 57850 120000 6 io_oeb[13]
port 69 nsew signal output
rlabel metal2 s 62118 119200 62174 120000 6 io_oeb[14]
port 70 nsew signal output
rlabel metal2 s 66350 119200 66406 120000 6 io_oeb[15]
port 71 nsew signal output
rlabel metal2 s 70674 119200 70730 120000 6 io_oeb[16]
port 72 nsew signal output
rlabel metal2 s 74998 119200 75054 120000 6 io_oeb[17]
port 73 nsew signal output
rlabel metal2 s 79230 119200 79286 120000 6 io_oeb[18]
port 74 nsew signal output
rlabel metal2 s 83554 119200 83610 120000 6 io_oeb[19]
port 75 nsew signal output
rlabel metal2 s 6366 119200 6422 120000 6 io_oeb[1]
port 76 nsew signal output
rlabel metal2 s 87786 119200 87842 120000 6 io_oeb[20]
port 77 nsew signal output
rlabel metal2 s 10690 119200 10746 120000 6 io_oeb[2]
port 78 nsew signal output
rlabel metal2 s 14922 119200 14978 120000 6 io_oeb[3]
port 79 nsew signal output
rlabel metal2 s 19246 119200 19302 120000 6 io_oeb[4]
port 80 nsew signal output
rlabel metal2 s 23478 119200 23534 120000 6 io_oeb[5]
port 81 nsew signal output
rlabel metal2 s 27802 119200 27858 120000 6 io_oeb[6]
port 82 nsew signal output
rlabel metal2 s 32126 119200 32182 120000 6 io_oeb[7]
port 83 nsew signal output
rlabel metal2 s 36358 119200 36414 120000 6 io_oeb[8]
port 84 nsew signal output
rlabel metal2 s 40682 119200 40738 120000 6 io_oeb[9]
port 85 nsew signal output
rlabel metal3 s 179200 14832 180000 14952 6 r
port 86 nsew signal output
rlabel metal3 s 0 17416 800 17536 6 rst
port 87 nsew signal input
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 88 nsew power input
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 88 nsew power input
rlabel metal4 s 65648 2128 65968 117552 6 vccd1
port 88 nsew power input
rlabel metal4 s 96368 2128 96688 117552 6 vccd1
port 88 nsew power input
rlabel metal4 s 127088 2128 127408 117552 6 vccd1
port 88 nsew power input
rlabel metal4 s 157808 2128 158128 117552 6 vccd1
port 88 nsew power input
rlabel metal3 s 0 24488 800 24608 6 vs
port 89 nsew signal output
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 90 nsew ground input
rlabel metal4 s 50288 2128 50608 117552 6 vssd1
port 90 nsew ground input
rlabel metal4 s 81008 2128 81328 117552 6 vssd1
port 90 nsew ground input
rlabel metal4 s 111728 2128 112048 117552 6 vssd1
port 90 nsew ground input
rlabel metal4 s 142448 2128 142768 117552 6 vssd1
port 90 nsew ground input
rlabel metal4 s 173168 2128 173488 117552 6 vssd1
port 90 nsew ground input
rlabel metal2 s 4066 0 4122 800 6 wbs_cyc_i
port 91 nsew signal input
rlabel metal2 s 12162 0 12218 800 6 wbs_stb_i
port 92 nsew signal input
rlabel metal3 s 0 31560 800 31680 6 web
port 93 nsew signal input
rlabel metal3 s 179200 24896 180000 25016 6 wmask0[0]
port 94 nsew signal input
rlabel metal2 s 113546 119200 113602 120000 6 wmask0[1]
port 95 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 180000 120000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 5981076
string GDS_FILE /home/fabio/chip_tutorial/upb_natalius_soc/openlane/natalius_soc/runs/natalius_soc/results/finishing/natalius_soc.magic.gds
string GDS_START 263090
<< end >>

